library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity g44_MAC_tb is
end g44_MAC_tb;
